module ALU_16_bit(
input wire [15:0] A,
input wire [15:0] B,
input wire [3:0] ALU_FUN,
input wire clk,
output reg [15:0] ALU_OUT,
output reg Carry_Flag,
output reg Arith_Flag,
output reg Logic_Flag,
output reg CMP_Flag,
output reg Shift_Flag
);

reg [15:0] ALU_OUT_Comb;

always @ (*)
 begin
  Arith_Flag = 0;
  Logic_Flag = 0;
  CMP_Flag = 0;
  Shift_Flag = 0;
	 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////	 
	 
  case (ALU_FUN)
    4'b0000: begin
	          {Carry_Flag, ALU_OUT_Comb} = A + B;
	          Arith_Flag = 1; 
			 end
 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	
	4'b0001: begin 
	          {Carry_Flag, ALU_OUT_Comb} = A - B;
	          Arith_Flag = 1;
 			 end
			 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	4'b0010: begin 
	          ALU_OUT_Comb = A * B;
	          Arith_Flag = 1; 
			 end
	
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	4'b0011: begin
	          if (B != 16'b0)
	           begin
			    ALU_OUT_Comb = A / B;
				Arith_Flag = 1;
			   end
			  else
			   begin
			    ALU_OUT_Comb = 16'b0;
				Arith_Flag = 1;
			   end
			 end
			   
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////			   

	4'b0100: begin 
	          ALU_OUT_Comb = A & B;
	          Logic_Flag = 1; 
			 end
			 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////			 
			 
	4'b0101: begin
	          ALU_OUT_Comb = A | B;
	          Logic_Flag = 1;
			 end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////			 
			 
	4'b0110: begin 
	          ALU_OUT_Comb = ~ (A & B);
	          Logic_Flag = 1;
			 end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////			 
			 
	4'b0111: begin
	          ALU_OUT_Comb = ~ (A | B);
	          Logic_Flag = 1;
			 end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	4'b1000: begin
	          ALU_OUT_Comb = A ^ B;
	          Logic_Flag = 1;
			 end
			 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////			 
			 
	4'b1001: begin 
	          ALU_OUT_Comb = ~ (A ^ B);
	          Logic_Flag = 1;
			 end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	4'b1010: begin
	          if (A == B)
	           begin
			    ALU_OUT_Comb = 16'b1;
				CMP_Flag = 1;
			   end
			  else
			   begin
			    ALU_OUT_Comb = 16'b0;
				CMP_Flag = 1;
			   end
			 end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	
	4'b1011: begin
	          if (A > B)
	           begin
			    ALU_OUT_Comb = 16'b10;
				CMP_Flag = 1;
			   end
			  else
			   begin
			    ALU_OUT_Comb = 16'b0;
				CMP_Flag = 1;
			   end
			 end
			 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	4'b1100: begin
	          if (A < B)
	           begin
			    ALU_OUT_Comb = 16'b11;
				CMP_Flag = 1;
			   end
			  else
			   begin
			    ALU_OUT_Comb = 16'b0;
				CMP_Flag = 1;
			   end
			 end
			 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
			
	4'b1101: begin 
	          ALU_OUT_Comb = A >> 1 ;
	          Shift_Flag = 1;
			 end
			 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	
	4'b1110: begin
           	  ALU_OUT_Comb = A << 1 ;
	          Shift_Flag = 1;
			 end
			 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////			 
			 
	default: ALU_OUT_Comb = 16'b0;
	
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	
  endcase
 end
 
always @ (posedge clk)
 begin
  ALU_OUT <= ALU_OUT_Comb;
 end 
	 
endmodule